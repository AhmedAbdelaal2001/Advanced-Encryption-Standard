//This module applies a substitution scheme to 1 byte of data.
//The substitution is as follows: compute the multiplicative inverse
//of the input data in the Galois field GF(2^8), and then apply the
//affine transformation shown in section 5.1.1.

module sBox(input[7:0] galoisField_byte,
				output reg[7:0] AffineTransformed_byte);
	//galoisField_byte: Input byte
	//AffineTransformed_byte: Output byte
	
	//Instead of implementing the extended Euclidean algorithm and the
	//affine transformation, the S-box will be used to compute the result.
	always @(*) 
	begin: substitution
		case(galoisField_byte)
			8'h00: AffineTransformed_byte=8'h63;
			8'h01: AffineTransformed_byte=8'h7c;
			8'h02: AffineTransformed_byte=8'h77;
			8'h03: AffineTransformed_byte=8'h7b;
			8'h04: AffineTransformed_byte=8'hf2;
			8'h05: AffineTransformed_byte=8'h6b;
			8'h06: AffineTransformed_byte=8'h6f;
			8'h07: AffineTransformed_byte=8'hc5;
			8'h08: AffineTransformed_byte=8'h30;
			8'h09: AffineTransformed_byte=8'h01;
			8'h0a: AffineTransformed_byte=8'h67;
			8'h0b: AffineTransformed_byte=8'h2b;
			8'h0c: AffineTransformed_byte=8'hfe;
			8'h0d: AffineTransformed_byte=8'hd7;
			8'h0e: AffineTransformed_byte=8'hab;
			8'h0f: AffineTransformed_byte=8'h76;
			8'h10: AffineTransformed_byte=8'hca;
			8'h11: AffineTransformed_byte=8'h82;
			8'h12: AffineTransformed_byte=8'hc9;
			8'h13: AffineTransformed_byte=8'h7d;
			8'h14: AffineTransformed_byte=8'hfa;
			8'h15: AffineTransformed_byte=8'h59;
			8'h16: AffineTransformed_byte=8'h47;
			8'h17: AffineTransformed_byte=8'hf0;
			8'h18: AffineTransformed_byte=8'had;
			8'h19: AffineTransformed_byte=8'hd4;
			8'h1a: AffineTransformed_byte=8'ha2;
			8'h1b: AffineTransformed_byte=8'haf;
			8'h1c: AffineTransformed_byte=8'h9c;
			8'h1d: AffineTransformed_byte=8'ha4;
			8'h1e: AffineTransformed_byte=8'h72;
			8'h1f: AffineTransformed_byte=8'hc0;
			8'h20: AffineTransformed_byte=8'hb7;
			8'h21: AffineTransformed_byte=8'hfd;
			8'h22: AffineTransformed_byte=8'h93;
			8'h23: AffineTransformed_byte=8'h26;
			8'h24: AffineTransformed_byte=8'h36;
			8'h25: AffineTransformed_byte=8'h3f;
			8'h26: AffineTransformed_byte=8'hf7;
			8'h27: AffineTransformed_byte=8'hcc;
			8'h28: AffineTransformed_byte=8'h34;
			8'h29: AffineTransformed_byte=8'ha5;
			8'h2a: AffineTransformed_byte=8'he5;
			8'h2b: AffineTransformed_byte=8'hf1;
			8'h2c: AffineTransformed_byte=8'h71;
			8'h2d: AffineTransformed_byte=8'hd8;
			8'h2e: AffineTransformed_byte=8'h31;
			8'h2f: AffineTransformed_byte=8'h15;
			8'h30: AffineTransformed_byte=8'h04;
			8'h31: AffineTransformed_byte=8'hc7;
			8'h32: AffineTransformed_byte=8'h23;
			8'h33: AffineTransformed_byte=8'hc3;
			8'h34: AffineTransformed_byte=8'h18;
			8'h35: AffineTransformed_byte=8'h96;
			8'h36: AffineTransformed_byte=8'h05;
			8'h37: AffineTransformed_byte=8'h9a;
			8'h38: AffineTransformed_byte=8'h07;
			8'h39: AffineTransformed_byte=8'h12;
			8'h3a: AffineTransformed_byte=8'h80;
			8'h3b: AffineTransformed_byte=8'he2;
			8'h3c: AffineTransformed_byte=8'heb;
			8'h3d: AffineTransformed_byte=8'h27;
			8'h3e: AffineTransformed_byte=8'hb2;
			8'h3f: AffineTransformed_byte=8'h75;
			8'h40: AffineTransformed_byte=8'h09;
			8'h41: AffineTransformed_byte=8'h83;
			8'h42: AffineTransformed_byte=8'h2c;
			8'h43: AffineTransformed_byte=8'h1a;
			8'h44: AffineTransformed_byte=8'h1b;
			8'h45: AffineTransformed_byte=8'h6e;
			8'h46: AffineTransformed_byte=8'h5a;
			8'h47: AffineTransformed_byte=8'ha0;
			8'h48: AffineTransformed_byte=8'h52;
			8'h49: AffineTransformed_byte=8'h3b;
			8'h4a: AffineTransformed_byte=8'hd6;
			8'h4b: AffineTransformed_byte=8'hb3;
			8'h4c: AffineTransformed_byte=8'h29;
			8'h4d: AffineTransformed_byte=8'he3;
			8'h4e: AffineTransformed_byte=8'h2f;
			8'h4f: AffineTransformed_byte=8'h84;
			8'h50: AffineTransformed_byte=8'h53;
			8'h51: AffineTransformed_byte=8'hd1;
			8'h52: AffineTransformed_byte=8'h00;
			8'h53: AffineTransformed_byte=8'hed;
			8'h54: AffineTransformed_byte=8'h20;
			8'h55: AffineTransformed_byte=8'hfc;
			8'h56: AffineTransformed_byte=8'hb1;
			8'h57: AffineTransformed_byte=8'h5b;
			8'h58: AffineTransformed_byte=8'h6a;
			8'h59: AffineTransformed_byte=8'hcb;
			8'h5a: AffineTransformed_byte=8'hbe;
			8'h5b: AffineTransformed_byte=8'h39;
			8'h5c: AffineTransformed_byte=8'h4a;
			8'h5d: AffineTransformed_byte=8'h4c;
			8'h5e: AffineTransformed_byte=8'h58;
			8'h5f: AffineTransformed_byte=8'hcf;
			8'h60: AffineTransformed_byte=8'hd0;
			8'h61: AffineTransformed_byte=8'hef;
			8'h62: AffineTransformed_byte=8'haa;
			8'h63: AffineTransformed_byte=8'hfb;
			8'h64: AffineTransformed_byte=8'h43;
			8'h65: AffineTransformed_byte=8'h4d;
			8'h66: AffineTransformed_byte=8'h33;
			8'h67: AffineTransformed_byte=8'h85;
			8'h68: AffineTransformed_byte=8'h45;
			8'h69: AffineTransformed_byte=8'hf9;
			8'h6a: AffineTransformed_byte=8'h02;
			8'h6b: AffineTransformed_byte=8'h7f;
			8'h6c: AffineTransformed_byte=8'h50;
			8'h6d: AffineTransformed_byte=8'h3c;
			8'h6e: AffineTransformed_byte=8'h9f;
			8'h6f: AffineTransformed_byte=8'ha8;
			8'h70: AffineTransformed_byte=8'h51;
			8'h71: AffineTransformed_byte=8'ha3;
			8'h72: AffineTransformed_byte=8'h40;
			8'h73: AffineTransformed_byte=8'h8f;
			8'h74: AffineTransformed_byte=8'h92;
			8'h75: AffineTransformed_byte=8'h9d;
			8'h76: AffineTransformed_byte=8'h38;
			8'h77: AffineTransformed_byte=8'hf5;
			8'h78: AffineTransformed_byte=8'hbc;
			8'h79: AffineTransformed_byte=8'hb6;
			8'h7a: AffineTransformed_byte=8'hda;
			8'h7b: AffineTransformed_byte=8'h21;
			8'h7c: AffineTransformed_byte=8'h10;
			8'h7d: AffineTransformed_byte=8'hff;
			8'h7e: AffineTransformed_byte=8'hf3;
			8'h7f: AffineTransformed_byte=8'hd2;
			8'h80: AffineTransformed_byte=8'hcd;
			8'h81: AffineTransformed_byte=8'h0c;
			8'h82: AffineTransformed_byte=8'h13;
			8'h83: AffineTransformed_byte=8'hec;
			8'h84: AffineTransformed_byte=8'h5f;
			8'h85: AffineTransformed_byte=8'h97;
			8'h86: AffineTransformed_byte=8'h44;
			8'h87: AffineTransformed_byte=8'h17;
			8'h88: AffineTransformed_byte=8'hc4;
			8'h89: AffineTransformed_byte=8'ha7;
			8'h8a: AffineTransformed_byte=8'h7e;
			8'h8b: AffineTransformed_byte=8'h3d;
			8'h8c: AffineTransformed_byte=8'h64;
			8'h8d: AffineTransformed_byte=8'h5d;
			8'h8e: AffineTransformed_byte=8'h19;
			8'h8f: AffineTransformed_byte=8'h73;
			8'h90: AffineTransformed_byte=8'h60;
			8'h91: AffineTransformed_byte=8'h81;
			8'h92: AffineTransformed_byte=8'h4f;
			8'h93: AffineTransformed_byte=8'hdc;
			8'h94: AffineTransformed_byte=8'h22;
			8'h95: AffineTransformed_byte=8'h2a;
			8'h96: AffineTransformed_byte=8'h90;
			8'h97: AffineTransformed_byte=8'h88;
			8'h98: AffineTransformed_byte=8'h46;
			8'h99: AffineTransformed_byte=8'hee;
			8'h9a: AffineTransformed_byte=8'hb8;
			8'h9b: AffineTransformed_byte=8'h14;
			8'h9c: AffineTransformed_byte=8'hde;
			8'h9d: AffineTransformed_byte=8'h5e;
			8'h9e: AffineTransformed_byte=8'h0b;
			8'h9f: AffineTransformed_byte=8'hdb;
			8'ha0: AffineTransformed_byte=8'he0;
			8'ha1: AffineTransformed_byte=8'h32;
			8'ha2: AffineTransformed_byte=8'h3a;
			8'ha3: AffineTransformed_byte=8'h0a;
			8'ha4: AffineTransformed_byte=8'h49;
			8'ha5: AffineTransformed_byte=8'h06;
			8'ha6: AffineTransformed_byte=8'h24;
			8'ha7: AffineTransformed_byte=8'h5c;
			8'ha8: AffineTransformed_byte=8'hc2;
			8'ha9: AffineTransformed_byte=8'hd3;
			8'haa: AffineTransformed_byte=8'hac;
			8'hab: AffineTransformed_byte=8'h62;
			8'hac: AffineTransformed_byte=8'h91;
			8'had: AffineTransformed_byte=8'h95;
			8'hae: AffineTransformed_byte=8'he4;
			8'haf: AffineTransformed_byte=8'h79;
			8'hb0: AffineTransformed_byte=8'he7;
			8'hb1: AffineTransformed_byte=8'hc8;
			8'hb2: AffineTransformed_byte=8'h37;
			8'hb3: AffineTransformed_byte=8'h6d;
			8'hb4: AffineTransformed_byte=8'h8d;
			8'hb5: AffineTransformed_byte=8'hd5;
			8'hb6: AffineTransformed_byte=8'h4e;
			8'hb7: AffineTransformed_byte=8'ha9;
			8'hb8: AffineTransformed_byte=8'h6c;
			8'hb9: AffineTransformed_byte=8'h56;
			8'hba: AffineTransformed_byte=8'hf4;
			8'hbb: AffineTransformed_byte=8'hea;
			8'hbc: AffineTransformed_byte=8'h65;
			8'hbd: AffineTransformed_byte=8'h7a;
			8'hbe: AffineTransformed_byte=8'hae;
			8'hbf: AffineTransformed_byte=8'h08;
			8'hc0: AffineTransformed_byte=8'hba;
			8'hc1: AffineTransformed_byte=8'h78;
			8'hc2: AffineTransformed_byte=8'h25;
			8'hc3: AffineTransformed_byte=8'h2e;
			8'hc4: AffineTransformed_byte=8'h1c;
			8'hc5: AffineTransformed_byte=8'ha6;
			8'hc6: AffineTransformed_byte=8'hb4;
			8'hc7: AffineTransformed_byte=8'hc6;
			8'hc8: AffineTransformed_byte=8'he8;
			8'hc9: AffineTransformed_byte=8'hdd;
			8'hca: AffineTransformed_byte=8'h74;
			8'hcb: AffineTransformed_byte=8'h1f;
			8'hcc: AffineTransformed_byte=8'h4b;
			8'hcd: AffineTransformed_byte=8'hbd;
			8'hce: AffineTransformed_byte=8'h8b;
			8'hcf: AffineTransformed_byte=8'h8a;
			8'hd0: AffineTransformed_byte=8'h70;
			8'hd1: AffineTransformed_byte=8'h3e;
			8'hd2: AffineTransformed_byte=8'hb5;
			8'hd3: AffineTransformed_byte=8'h66;
			8'hd4: AffineTransformed_byte=8'h48;
			8'hd5: AffineTransformed_byte=8'h03;
			8'hd6: AffineTransformed_byte=8'hf6;
			8'hd7: AffineTransformed_byte=8'h0e;
			8'hd8: AffineTransformed_byte=8'h61;
			8'hd9: AffineTransformed_byte=8'h35;
			8'hda: AffineTransformed_byte=8'h57;
			8'hdb: AffineTransformed_byte=8'hb9;
			8'hdc: AffineTransformed_byte=8'h86;
			8'hdd: AffineTransformed_byte=8'hc1;
			8'hde: AffineTransformed_byte=8'h1d;
			8'hdf: AffineTransformed_byte=8'h9e;
			8'he0: AffineTransformed_byte=8'he1;
			8'he1: AffineTransformed_byte=8'hf8;
			8'he2: AffineTransformed_byte=8'h98;
			8'he3: AffineTransformed_byte=8'h11;
			8'he4: AffineTransformed_byte=8'h69;
			8'he5: AffineTransformed_byte=8'hd9;
			8'he6: AffineTransformed_byte=8'h8e;
			8'he7: AffineTransformed_byte=8'h94;
			8'he8: AffineTransformed_byte=8'h9b;
			8'he9: AffineTransformed_byte=8'h1e;
			8'hea: AffineTransformed_byte=8'h87;
			8'heb: AffineTransformed_byte=8'he9;
			8'hec: AffineTransformed_byte=8'hce;
			8'hed: AffineTransformed_byte=8'h55;
			8'hee: AffineTransformed_byte=8'h28;
			8'hef: AffineTransformed_byte=8'hdf;
			8'hf0: AffineTransformed_byte=8'h8c;
			8'hf1: AffineTransformed_byte=8'ha1;
			8'hf2: AffineTransformed_byte=8'h89;
			8'hf3: AffineTransformed_byte=8'h0d;
			8'hf4: AffineTransformed_byte=8'hbf;
			8'hf5: AffineTransformed_byte=8'he6;
			8'hf6: AffineTransformed_byte=8'h42;
			8'hf7: AffineTransformed_byte=8'h68;
			8'hf8: AffineTransformed_byte=8'h41;
			8'hf9: AffineTransformed_byte=8'h99;
			8'hfa: AffineTransformed_byte=8'h2d;
			8'hfb: AffineTransformed_byte=8'h0f;
			8'hfc: AffineTransformed_byte=8'hb0;
			8'hfd: AffineTransformed_byte=8'h54;
			8'hfe: AffineTransformed_byte=8'hbb;
			8'hff: AffineTransformed_byte=8'h16;
		endcase
	end
endmodule
